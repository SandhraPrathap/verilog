// Code your design here
module and_2_datafl(input A,input B, output Y);
assign Y = A & B; 
endmodule 