module and_2_str(input A, input B, output Y);

  and and1 (Y, A, B);
  endmodule